`include "D:/uvm_proj/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqNNNN.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqNNN.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqNNNNQ.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqNDN.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqNDNN.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqDNND.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqDNN.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqDNNN.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqNDND.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqQ.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqNNNND.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqNNNNN.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqNNDQ.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqDDN.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqNNND.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqNDQ.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqND.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqNDNQ.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqDND.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqDDD.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqNN.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqNNNQ.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqNQ.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqNNQ.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqN.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqDD.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqNND.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqNNDN.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqDDQ.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqDNQ.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqD.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqDNNQ.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqDN.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqDQ.sv"
