// ----------- ---------- candy_vending_seqNNNND.sv	candy_vending_seqNNNND	seqNNNND_tx  ----------- ---------- 
// ----------- ---------- D:/uvm_proj/acvm_new/candy_vending_DV/cv_agent/cv_sequences/candy_vending_seqNNNND.sv ----------- ---------- 
class candy_vending_seqNNNND extends uvm_sequence#(candy_vending_seq_item);
	`uvm_object_utils(candy_vending_seqNNNND)


	function new(string name = "");
		super.new(name);
	endfunction

	task body();

		set_response_queue_error_report_disabled(1);

		repeat (10) begin

			candy_vending_seq_item seqNNNND_tx;
			seqNNNND_tx = new ("seqNNNND_tx");

			seqNNNND_tx = candy_vending_seq_item::type_id::create("seqNNNND_tx");
			start_item(seqNNNND_tx);


			// randomize the sequence or assign values for respective seq items
			//seqNNNND_tx.coins = {N,N,N,N,D};
			//seqNNNND_tx.cancel = 0;


			// Trying to randomize dynamic array with inline constraint, results in error

			void'(seqNNNND_tx.randomize() with {coin_cnt == 5; cost== 30 ; cancel == 0 ;}); // inline type

			`uvm_info("SEQUENCE_NNNND",$sformatf ("no of coins %0d", seqNNNND_tx.coins.size()),UVM_LOW);
	
				`uvm_info("SEQUENCE_NNNND",$sformatf ("coins are %0s,%0s,%0s,%0s,%0s !",seqNNNND_tx.coins[4],seqNNNND_tx.coins[3],seqNNNND_tx.coins[2],seqNNNND_tx.coins[1],seqNNNND_tx.coins[0]),UVM_LOW);

				`uvm_info(get_type_name(),seq20_tx.convert2string(),UVM_LOW);
			finish_item(seqNNNND_tx);
		end
	endtask

endclass


//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


