`include "D:/uvm_proj/candy_vending_DV/cv_tests/candy_vending_testcaseNNNN.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_tests/candy_vending_testcaseNNN.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_tests/candy_vending_testcaseNNNNQ.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_tests/candy_vending_testcaseNDN.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_tests/candy_vending_testcaseNDNN.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_tests/candy_vending_testcaseDNND.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_tests/candy_vending_testcaseDNN.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_tests/candy_vending_testcaseDNNN.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_tests/candy_vending_testcaseNDND.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_tests/candy_vending_testcaseQ.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_tests/candy_vending_testcaseNNNND.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_tests/candy_vending_testcaseNNNNN.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_tests/candy_vending_testcaseNNDQ.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_tests/candy_vending_testcaseDDN.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_tests/candy_vending_testcaseNNND.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_tests/candy_vending_testcaseNDQ.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_tests/candy_vending_testcaseND.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_tests/candy_vending_testcaseNDNQ.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_tests/candy_vending_testcaseDND.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_tests/candy_vending_testcaseDDD.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_tests/candy_vending_testcaseNN.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_tests/candy_vending_testcaseNNNQ.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_tests/candy_vending_testcaseNQ.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_tests/candy_vending_testcaseNNQ.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_tests/candy_vending_testcaseN.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_tests/candy_vending_testcaseDD.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_tests/candy_vending_testcaseNND.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_tests/candy_vending_testcaseNNDN.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_tests/candy_vending_testcaseDDQ.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_tests/candy_vending_testcaseDNQ.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_tests/candy_vending_testcaseD.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_tests/candy_vending_testcaseDNNQ.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_tests/candy_vending_testcaseDN.sv"
`include "D:/uvm_proj/candy_vending_DV/cv_tests/candy_vending_testcaseDQ.sv"
